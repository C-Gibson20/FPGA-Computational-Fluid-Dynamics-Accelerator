module SolverDMA_top (
    ports
);
    
endmodule