module image_thing2 (
    input wire [31:0] din,
    input wire [31:0] addr,
    input wire clk
);


    

endmodule