`ifndef DEF
`define DEF

`define DATA_WIDTH 16
`define HEIGHT 300
`define WIDTH 100
`define DEPTH (HEIGHT*WIDTH)
`define ADDRESS_WIDTH ($clog2(DEPTH))

`endif
