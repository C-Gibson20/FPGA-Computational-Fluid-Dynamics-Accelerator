`include "def.sv"

module LBMSolver (
    input logic clk,
    input logic rst, 
    input logic en
);

logic [`DATA_WIDTH-1:0] c0_data_in, c0_data_out;
logic c0_mem_write;
logic [`ADDRESS_WIDTH-1:0] c0_write_address,c0_read_address;

logic [`DATA_WIDTH-1:0] cn_data_in , cn_data_out;
logic cn_mem_write;
logic [`ADDRESS_WIDTH-1:0] cn_write_address, cn_read_address;

logic [`DATA_WIDTH-1:0] cne_data_in, cne_data_out;
logic cne_mem_write;
logic [`ADDRESS_WIDTH-1:0] cne_write_address,cne_read_address;

logic [`DATA_WIDTH-1:0] ce_data_in ,ce_data_out;
logic ce_mem_write;
logic [`ADDRESS_WIDTH-1:0] ce_write_address, ce_read_address;

logic [`DATA_WIDTH-1:0] cse_data_in , cse_data_out;
logic cse_mem_write;
logic [`ADDRESS_WIDTH-1:0] cse_write_address, cse_read_address;

logic [`DATA_WIDTH-1:0] cs_data_in, cs_data_out;
logic cs_mem_write;
logic [`ADDRESS_WIDTH-1:0] cs_write_address, cs_read_address;

logic [`DATA_WIDTH-1:0] csw_data_in, csw_data_out;
logic csw_mem_write;
logic [`ADDRESS_WIDTH-1:0] csw_write_address, csw_read_address;

logic [`DATA_WIDTH-1:0] cw_data_in, cw_data_out;
logic cw_mem_write;
logic [`ADDRESS_WIDTH-1:0] cw_write_address, cw_read_address;

logic [`DATA_WIDTH-1:0] cnw_data_in, cnw_data_out;
logic cnw_mem_write;
logic [`ADDRESS_WIDTH-1:0] cnw_write_address, cnw_read_address;

//Stores the 9 directions in their own RAM, I can't make each cell it's own block of memory, so instead I've decided to split the memory by direction
RAM C0(
    .read_address(c0_read_address),
    .write_address(c0_write_address),
    .data_in(c0_data_in),
    .clk(clk),
    .mem_write(c0_mem_write),
    .data_out(c0_data_out)
);

RAM CN(
    .read_address(cn_read_address),
    .write_address(cn_write_address),
    .data_in(cn_data_in),
    .clk(clk),
    .mem_write(cn_mem_write),
    .data_out(cn_data_out)
);

RAM CNE(
    .read_address(cne_read_address),
    .write_address(cne_write_address),
    .data_in(cne_data_in),
    .clk(clk),
    .mem_write(cne_mem_write),
    .data_out(cne_data_out)
);

RAM CE(
    .read_address(ce_read_address),
    .write_address(ce_write_address),
    .data_in(ce_data_in),
    .clk(clk),
    .mem_write(ce_mem_write),
    .data_out(ce_data_out)
);

RAM CSE(
    .read_address(cse_read_address),
    .write_address(cse_write_address),
    .data_in(cse_data_in),
    .clk(clk),
    .mem_write(cse_mem_write),
    .data_out(cse_data_out)
);

RAM CS(
    .read_address(cs_read_address),
    .write_address(cs_write_address),
    .data_in(cs_data_in),
    .clk(clk),
    .mem_write(cs_mem_write),
    .data_out(cs_data_out)
);

RAM CSW(
    .read_address(csw_read_address),
    .write_address(csw_write_address),
    .data_in(csw_data_in),
    .clk(clk),
    .mem_write(csw_mem_write),
    .data_out(csw_data_out)
);

RAM CW(
    .read_address(cw_read_address),
    .write_address(cw_write_address),
    .data_in(cw_data_in),
    .clk(clk),
    .mem_write(cw_mem_write),
    .data_out(cw_data_out)
);

RAM CNW(
    .read_address(cnw_read_address),
    .write_address(cnw_write_address),
    .data_in(cnw_data_in),
    .clk(clk),
    .mem_write(cnw_mem_write),
    .data_out(cnw_data_out)
);


endmodule
