module top #(
    parameters
) (
    ports
);
    
endmodule